--
-- VHDL Architecture ece411.X3b.untitled
--
-- Created:
--          by - tischer1.ews (evrt-252-20.ews.illinois.edu)
--          at - 18:58:16 11/13/12
--
-- using Mentor Graphics HDL Designer(TM) 2005.3 (Build 75)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY X3b IS
   PORT( 
      x3out : OUT    LC3b_reg
   );

-- Declarations

END X3b ;

--
ARCHITECTURE untitled OF X3b IS
BEGIN
  x3out <= "XXX";
END ARCHITECTURE untitled;

