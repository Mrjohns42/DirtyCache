--
-- VHDL Architecture ece411.RegFile.untitled
--
-- Created:
--          by - hcander2.ews (linux7.ews.illinois.edu)
--          at - 02:03:28 09/05/12
--
-- using Mentor Graphics HDL Designer(TM) 2005.3 (Build 75)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY RegFile IS
   PORT( 
      Dest     : IN     LC3b_reg;
      reset_l  : IN     std_logic;
      Input    : IN     LC3b_word;
      RegWrite : IN     std_logic;
      SrcB     : IN     LC3b_reg;
      SrcA     : IN     LC3b_reg;
      clk      : IN     std_logic;
      RFA      : OUT    LC3b_word;
      RFB      : OUT    LC3b_word
   );

-- Declarations

END RegFile ;

--
ARCHITECTURE untitled OF RegFile IS
TYPE RAMMEMORY IS ARRAY (7 DOWNTO 0) OF LC3b_word;
SIGNAL RAM : RAMMEMORY;
BEGIN
  -------------------------------------------------------------------
  VHDL_REGFILE_READ : PROCESS (RAM, SrcA, SrcB)
  -------------------------------------------------------------------
  VARIABLE RADDR1 : INTEGER RANGE 0 TO 7;
  VARIABLE RADDR2 : INTEGER RANGE 0 TO 7;
  BEGIN
    --READ FROM REGFILE, THE OUTPUTS ARE VALID AFTER REGFILE_READ DELAY.
    RADDR1 := TO_INTEGER(UNSIGNED('0' & SrcA));
    RADDR2 := TO_INTEGER(UNSIGNED('0' & SrcB));
    RFA <= RAM(RADDR1) AFTER DELAY_REGFILE_READ;
    RFB <= RAM(RADDR2) AFTER DELAY_REGFILE_READ;
  END PROCESS VHDL_REGFILE_READ;
  -------------------------------------------------------------------
  VHDL_REGFILE_WRITE: PROCESS(clk, Input, RegWrite, Dest, reset_l)
  -------------------------------------------------------------------
  VARIABLE WADDR : INTEGER RANGE 0 TO 7;
  BEGIN
    -- ON RESET, CLEAR THE REGISTER FILE CONTENTS
    IF (reset_l = '0') THEN
      RAM(0) <= "0000000000000000";
      RAM(1) <= "0000000000000000";
      RAM(2) <= "0000000000000000";
      RAM(3) <= "0000000000000000";
      RAM(4) <= "0000000000000000";
      RAM(5) <= "0000000000000000";
      RAM(6) <= "0000000000000000";
      RAM(7) <= "0000000000000000";
    END IF;
    -- WRITE VALUE TO REGISTER FILE ON RISING EDGE OF CLOCK IF REGWRITE ACTIVE
    -- NOW FALLING EDGE FOR FORWARDING
    WADDR := TO_INTEGER(UNSIGNED('0' & Dest));
    IF (CLK'EVENT AND (clk = '0') AND (CLK'LAST_VALUE = '1')) THEN
      IF (RegWrite = '1') THEN
        RAM(WADDR) <= Input;
      END IF;
    END IF;
  END PROCESS VHDL_REGFILE_WRITE;
END ARCHITECTURE untitled;

